`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date:    21:01:40 05/22/2019
// Design Name:
// Module Name:    id_exe_register
// Project Name:
// Target Devices:
// Tool versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
module id_exe_register(clk,clrn,
                       lock_write, // stall 锁住写信号，消除指令的影响
                       id_wreg,id_m2reg,id_wmem,id_aluc,id_aluimm,id_a,id_b,id_imm,id_rn,id_shift,id_wz,
                       exe_wreg,exe_m2reg,exe_wmem,exe_aluc,exe_aluimm,exe_a,exe_b,exe_imm,exe_rn,exe_shift,exe_wz
                      );
input [31:0] id_a,id_b,id_imm;
input [4:0] id_rn;
input [2:0] id_aluc;
input id_wreg,id_m2reg,id_wmem,id_aluimm,id_shift,id_wz;
input clk,clrn, lock_write;

output reg [31:0] exe_a,exe_b,exe_imm;
output reg [4:0] exe_rn;
output reg [2:0] exe_aluc;
output reg exe_wreg,exe_m2reg,exe_wmem,exe_aluimm,exe_shift,exe_wz;

//请在下方补充代码以完成流水线寄存器
//////////////////////////////////////////////////////////////////////////////

always @(posedge clk or negedge clrn) begin
    if (clrn == 0) begin
        exe_a <= 0;
        exe_b <= 0;
        exe_imm <= 0;
        exe_rn <= 0;
        exe_aluc <= 0;

        exe_wreg <= 0;
        exe_m2reg <= 0;
        exe_wmem <= 0;
        exe_aluimm <= 0;
        exe_shift <= 0;
        exe_wz <= 0;
    end
    else if (lock_write) begin
        exe_wreg <= 0;
        exe_wz <= 0;
        exe_wmem <= 0;
    end
    else begin
        exe_a <= id_a;
        exe_b <= id_b;
        exe_imm <= id_imm;
        exe_rn <= id_rn;
        exe_aluc <= id_aluc;

        exe_wreg <= id_wreg;
        exe_wz <= id_wz;
        exe_wmem <= id_wmem;

        exe_m2reg <= id_m2reg;
        exe_aluimm <= id_aluimm;
        exe_shift <= id_shift;
    end
end

endmodule
